library ieee;
use ieee.std_logic_1164.all;

architecture beh of cnt_to_vga is
begin

end architecture beh;
